library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity testbench is
end testbench;

architecture tb of testbench is

signal A,B,R:bit_vector(15 downto 0);
signal P0,P1,C0,Z0:bit;

component ALU is
   Port( I0: in bit_vector(15 downto 0);
		I1: in bit_vector(15 downto 0);
		
		S0: in bit; --Control (select) Inputs
		S1: in bit;
		
		A: out bit_vector(15 downto 0);  --Output vector
		C: out bit;  --Carry
		Z: out bit);  --Zero bit
end component;


begin 
dut_instance:ALU
port map(I0=>A,I1=>B,S0=>P0, S1=>P1, A=>R,C=>C0,Z=>Z0);

process
begin

P0 <= '0';
P1 <= '0';
A<="0010001011111010";
B<="0010001011111010";

wait for 5 ns;
assert (R="0100010111110100" and C0='0' and Z0='1') report "testbench 1 is not ok";
wait for 5 ns;


P0 <= '0';
P1 <= '1';
A<="0010001011111010";
B<="0010001011111010";

wait for 5 ns;
assert (R="0000000000000000" and C0='0' and Z0='1') report "testbench 2 is not ok";
wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="0010001011111010";
B<="0010001011111010";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="0010001011111010";
B<="0010001011111010";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="0111000100000111";
B<="0101111101011101";

wait for 5 ns;


P0 <= '0';
P1 <= '1';
A<="0111000100000111";
B<="0101111101011101";

wait for 5 ns;


P0 <= '1';
P1 <= '0';
A<="0111000100000111";
B<="0101111101011101";

wait for 5 ns;


P0 <= '1';
P1 <= '1';
A<="0111000100000111";
B<="0101111101011101";

wait for 5 ns;


P0 <= '0';
P1 <= '0';
A<="0110001000001111";
B<="1111010011111100";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="0110001000001111";
B<="1111010011111100";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="0110001000001111";
B<="1111010011111100";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="0110001000001111";
B<="1111010011111100";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="0000011010010111";
B<="1110000100101010";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="0000011010010111";
B<="1110000100101010";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="0000011010010111";
B<="1110000100101010";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="0000011010010111";
B<="1110000100101010";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1010000101111011";
B<="0010001000110101";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1010000101111011";
B<="0010001000110101";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="1010000101111011";
B<="0010001000110101";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1010000101111011";
B<="0010001000110101";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1101000111111010";
B<="0101111011101000";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1101000111111010";
B<="0101111011101000";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="1101000111111010";
B<="0101111011101000";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1101000111111010";
B<="0101111011101000";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1100000011100000";
B<="1101010011111101";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1100000011100000";
B<="1101010011111101";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="1100000011100000";
B<="1101010011111101";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1100000011100000";
B<="1101010011111101";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1000111110010001";
B<="1000101000100111";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1000111110010001";
B<="1000101000100111";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="1000111110010001";
B<="1000101000100111";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1000111110010001";
B<="1000101000100111";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="0000000000000000";
B<="0000000000000000";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="0000000000000000";
B<="0000000000000000";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="0000000000000000";
B<="0000000000000000";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="0000000000000000";
B<="0000000000000000";

wait for 5 ns;


P0 <= '0';
P1 <= '0';
A<="0000000000000000";
B<="1111111111111111";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="0000000000000000";
B<="1111111111111111";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="0000000000000000";
B<="1111111111111111";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="0000000000000000";
B<="1111111111111111";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1111111111111111";
B<="0000000000000000";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1111111111111111";
B<="0000000000000000";

wait for 5 ns;
P0 <= '1';
P1 <= '0';
A<="1111111111111111";
B<="0000000000000000";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1111111111111111";
B<="0000000000000000";

wait for 5 ns;

P0 <= '0';
P1 <= '0';
A<="1111111111111111";
B<="1111111111111111";

wait for 5 ns;

P0 <= '0';
P1 <= '1';
A<="1111111111111111";
B<="1111111111111111";

wait for 5 ns;

P0 <= '1';
P1 <= '0';
A<="1111111111111111";
B<="1111111111111111";

wait for 5 ns;

P0 <= '1';
P1 <= '1';
A<="1111111111111111";
B<="1111111111111111";

wait for 5 ns;

end process;
end tb;